// ==========================================================
// Data Assembler
// ==========================================================
module data_assembler (
    input [511:0] lidar_data,
    input lidar_valid,
    input [3071:0] camera_data,
    input camera_valid,
    input [127:0] radar_data,
    input radar_valid,
    input [63:0] imu_data,
    input imu_valid,
    output logic [3839:0] fused_data,
    output logic valid
);

    always_comb begin
        valid = lidar_valid & camera_valid & radar_valid & imu_valid;
        if (valid) {
            fused_data[3839:3328] = lidar_data;
            fused_data[3327:256] = camera_data;
            fused_data[255:128] = radar_data;
            fused_data[127:64] = imu_data;
        } else {
            fused_data = '0;
        }
    end
endmodule

// ==========================================================
// Interpolation Calculator (fixed-point)
// ==========================================================
module interpolation_calculator #(
    parameter DATA_WIDTH = 512
)(
    input clk,
    input rst_n,
    input [63:0] t_common,
    input [DATA_WIDTH+63:0] packet1,
    input [DATA_WIDTH+63:0] packet2,
    input start,
    output logic [DATA_WIDTH-1:0] interpolated_data,
    output logic valid,
    output logic error
);

    logic [63:0] ts1, ts2;
    logic [DATA_WIDTH-1:0] data1, data2;
    logic [31:0] ratio;
    
    assign ts1 = packet1[DATA_WIDTH +: 64];
    assign ts2 = packet2[DATA_WIDTH +: 64];
    assign data1 = packet1[0 +: DATA_WIDTH];
    assign data2 = packet2[0 +: DATA_WIDTH];

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            interpolated_data <= 0;
            valid <= 0;
            error <= 0;
        end else if (start) begin
            valid <= 0;
            error <= 0;
            if (ts1 == t_common) begin
                interpolated_data <= data1;
                valid <= 1;
            end else if (ts2 == t_common) begin
                interpolated_data <= data2;
                valid <= 1;
            end else if (ts1 > t_common || ts2 < t_common) begin
                error <= 1;
            end else if (ts1 == ts2) begin
                interpolated_data <= data1;
                valid <= 1;
                error <= (ts1 != t_common);
            end else begin
                ratio = ((t_common - ts1) << 16) / (ts2 - ts1);
                for (int i = 0; i < DATA_WIDTH/32; i++) begin
                    logic [31:0] val1 = data1[i*32 +: 32];
                    logic [31:0] val2 = data2[i*32 +:32];
                    logic signed [31:0] delta = val2 - val1;
                    interpolated_data[i*32 +: 32] = val1 + ((delta * ratio) >> 16);
                end
                valid <= 1;
            end
        end else begin
            valid <= 0;
        end
    end
endmodule

// ==========================================================
// Matcher Unit (with binary search)
// ==========================================================
module matcher_unit #(
    parameter DATA_WIDTH = 512,
    parameter BUFFER_DEPTH = 16
)(
    input clk,
    input rst_n,
    input [63:0] t_common,
    input start,
    output logic done,
    output logic error,
    output logic [DATA_WIDTH+63:0] packet1,
    output logic [DATA_WIDTH+63:0] packet2,
    input [DATA_WIDTH+63:0] fifo_dout,
    input fifo_empty,
    output logic fifo_rd_en,
    input [ADDR_WIDTH:0] fifo_count
);

    localparam ADDR_WIDTH = $clog2(BUFFER_DEPTH);
    
    typedef enum {
        IDLE,
        INIT_SEARCH,
        BINARY_SEARCH,
        READ_SAMPLES,
        OUTPUT_DATA,
        ERROR_STATE
    } state_t;

    state_t state;
    logic [ADDR_WIDTH-1:0] low_ptr, high_ptr, mid_ptr;
    logic [63:0] mid_ts;
    logic found;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            done <= 0;
            error <= 0;
            fifo_rd_en <= 0;
            packet1 <= 0;
            packet2 <= 0;
        end else begin
            case (state)
                IDLE: begin
                    if (start && fifo_count >= 2) begin
                        state <= INIT_SEARCH;
                        low_ptr <= 0;
                        high_ptr <= fifo_count - 1;
                        found <= 0;
                    end else if (start) begin
                        state <= ERROR_STATE;
                    end
                end
                INIT_SEARCH: begin
                    state <= BINARY_SEARCH;
                end
                BINARY_SEARCH: begin
                    if (low_ptr <= high_ptr) begin
                        mid_ptr = low_ptr + ((high_ptr - low_ptr) >> 1);
                        fifo_rd_en <= 1;
                        state <= READ_MID;
                    end else begin
                        state <= ERROR_STATE;
                    end
                end
                READ_MID: begin
                    fifo_rd_en <= 0;
                    mid_ts <= fifo_dout[DATA_WIDTH +: 64];
                    if (mid_ts == t_common) begin
                        packet1 <= fifo_dout;
                        packet2 <= fifo_dout;
                        found <= 1;
                        state <= OUTPUT_DATA;
                    end else if (mid_ts < t_common) begin
                        low_ptr <= mid_ptr + 1;
                        state <= BINARY_SEARCH;
                    end else begin
                        high_ptr <= mid_ptr - 1;
                        state <= BINARY_SEARCH;
                    end
                end
                OUTPUT_DATA: begin
                    if (found) begin
                        done <= 1;
                        state <= IDLE;
                    end else begin
                        fifo_rd_en <= 1;
                        state <= READ_SAMPLES;
                    end
                end
                READ_SAMPLES: begin
                    packet1 <= fifo_dout;
                    fifo_rd_en <= 1;
                    packet2 <= fifo_dout;
                    state <= OUTPUT_DATA;
                end
                ERROR_STATE: begin
                    error <= 1;
                    done <= 1;
                    state <= IDLE;
                end
            endcase
        end
    end
endmodule


// ==========================================================
// Sensor Data Buffer (FIFO with timestamp)
// ==========================================================
module sensor_data_buffer #(
    parameter DATA_WIDTH = 512,
    parameter BUFFER_DEPTH = 16,
    parameter ADDR_WIDTH = $clog2(BUFFER_DEPTH)
)(
    input clk,
    input rst_n,
    input wr_en,
    input [DATA_WIDTH+63:0] din,  // {data, timestamp}
    input rd_en,
    output logic [DATA_WIDTH+63:0] dout,
    output logic full,
    output logic empty,
    output logic [ADDR_WIDTH:0] count
);

    logic [DATA_WIDTH+63:0] mem [0:BUFFER_DEPTH-1];
    logic [ADDR_WIDTH-1:0] wr_ptr, rd_ptr;
    logic [ADDR_WIDTH:0] item_count;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            wr_ptr <= 0;
            rd_ptr <= 0;
            item_count <= 0;
            empty <= 1;
            full <= 0;
            for (int i = 0; i < BUFFER_DEPTH; i++) mem[i] <= 0;
        end else begin
            if (wr_en && !full) begin
                mem[wr_ptr] <= din;
                wr_ptr <= (wr_ptr == BUFFER_DEPTH-1) ? 0 : wr_ptr + 1;
                item_count <= item_count + 1;
            end
            if (rd_en && !empty) begin
                dout <= mem[rd_ptr];
                rd_ptr <= (rd_ptr == BUFFER_DEPTH-1) ? 0 : rd_ptr + 1;
                item_count <= item_count - 1;
            end
            empty <= (item_count == 0);
            full <= (item_count == BUFFER_DEPTH);
        end
    end

    assign count = item_count;
endmodule

// ==========================================================
// Time Reference Module
// ==========================================================
module time_reference (
    input clk,
    input rst_n,
    input sync_signal,
    output logic [63:0] t_common
);

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            t_common <= 0;
        end else if (sync_signal) begin
            t_common <= t_common + 1;
        end
    end
endmodule


// ==========================================================
// Timestamp Extractor
// ==========================================================
module timestamp_extractor #(
    parameter DATA_WIDTH = 512
)(
    input [DATA_WIDTH+63:0] data_in,
    output logic [63:0] timestamp,
    output logic [DATA_WIDTH-1:0] sensor_data
);
    assign timestamp = data_in[DATA_WIDTH +: 64];
    assign sensor_data = data_in[0 +: DATA_WIDTH];
endmodule


// ==========================================================
// Top-Level Temporal Alignment
// ==========================================================
module temporal_alignment (
    input clk,
    input rst_n,
    input sync_signal,
    input [575:0] lidar_din,
    input lidar_wr_en,
    input [3135:0] camera_din,
    input camera_wr_en,
    input [191:0] radar_din,
    input radar_wr_en,
    input [127:0] imu_din,
    input imu_wr_en,
    output logic [3839:0] fused_data,
    output logic valid,
    output logic error
);

    logic [63:0] t_common;
    time_reference time_ref (
        .clk(clk),
        .rst_n(rst_n),
        .sync_signal(sync_signal),
        .t_common(t_common)
    );

    logic [575:0] lidar_dout;
    logic [3135:0] camera_dout;
    logic [191:0] radar_dout;
    logic [127:0] imu_dout;
    
    logic lidar_empty, camera_empty, radar_empty, imu_empty;
    logic lidar_full, camera_full, radar_full, imu_full;
    logic lidar_rd_en, camera_rd_en, radar_rd_en, imu_rd_en;
    
    logic [3:0] lidar_count, camera_count, radar_count, imu_count;

    sensor_data_buffer #(
        .DATA_WIDTH(512),
        .BUFFER_DEPTH(16)
    ) lidar_buffer (
        .clk(clk),
        .rst_n(rst_n),
        .wr_en(lidar_wr_en),
        .din(lidar_din),
        .rd_en(lidar_rd_en),
        .dout(lidar_dout),
        .full(lidar_full),
        .empty(lidar_empty),
        .count(lidar_count)
    );

    sensor_data_buffer #(
        .DATA_WIDTH(3072),
        .BUFFER_DEPTH(16)
    ) camera_buffer (
        .clk(clk),
        .rst_n(rst_n),
        .wr_en(camera_wr_en),
        .din(camera_din),
        .rd_en(camera_rd_en),
        .dout(camera_dout),
        .full(camera_full),
        .empty(camera_empty),
        .count(camera_count)
    );

    sensor_data_buffer #(
        .DATA_WIDTH(128),
        .BUFFER_DEPTH(16)
    ) radar_buffer (
        .clk(clk),
        .rst_n(rst_n),
        .wr_en(radar_wr_en),
        .din(radar_din),
        .rd_en(radar_rd_en),
        .dout(radar_dout),
        .full(radar_full),
        .empty(radar_empty),
        .count(radar_count)
    );

    sensor_data_buffer #(
        .DATA_WIDTH(64),
        .BUFFER_DEPTH(16)
    ) imu_buffer (
        .clk(clk),
        .rst_n(rst_n),
        .wr_en(imu_wr_en),
        .din(imu_din),
        .rd_en(imu_rd_en),
        .dout(imu_dout),
        .full(imu_full),
        .empty(imu_empty),
        .count(imu_count)
    );

    logic [575:0] lidar_packet1, lidar_packet2;
    logic [3135:0] camera_packet1, camera_packet2;
    logic [191:0] radar_packet1, radar_packet2;
    logic [127:0] imu_packet1, imu_packet2;
    
    logic lidar_matcher_done, camera_matcher_done, radar_matcher_done, imu_matcher_done;
    logic lidar_matcher_error, camera_matcher_error, radar_matcher_error, imu_matcher_error;

    matcher_unit #(
        .DATA_WIDTH(512),
        .BUFFER_DEPTH(16)
    ) lidar_matcher (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .start(sync_signal),
        .done(lidar_matcher_done),
        .error(lidar_matcher_error),
        .packet1(lidar_packet1),
        .packet2(lidar_packet2),
        .fifo_dout(lidar_dout),
        .fifo_empty(lidar_empty),
        .fifo_rd_en(lidar_rd_en),
        .fifo_count(lidar_count)
    );

    matcher_unit #(
        .DATA_WIDTH(3072),
        .BUFFER_DEPTH(16)
    ) camera_matcher (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .start(sync_signal),
        .done(camera_matcher_done),
        .error(camera_matcher_error),
        .packet1(camera_packet1),
        .packet2(camera_packet2),
        .fifo_dout(camera_dout),
        .fifo_empty(camera_empty),
        .fifo_rd_en(camera_rd_en),
        .fifo_count(camera_count)
    );

    matcher_unit #(
        .DATA_WIDTH(128),
        .BUFFER_DEPTH(16)
    ) radar_matcher (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .start(sync_signal),
        .done(radar_matcher_done),
        .error(radar_matcher_error),
        .packet1(radar_packet1),
        .packet2(radar_packet2),
        .fifo_dout(radar_dout),
        .fifo_empty(radar_empty),
        .fifo_rd_en(radar_rd_en),
        .fifo_count(radar_count)
    );

    matcher_unit #(
        .DATA_WIDTH(64),
        .BUFFER_DEPTH(16)
    ) imu_matcher (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .start(sync_signal),
        .done(imu_matcher_done),
        .error(imu_matcher_error),
        .packet1(imu_packet1),
        .packet2(imu_packet2),
        .fifo_dout(imu_dout),
        .fifo_empty(imu_empty),
        .fifo_rd_en(imu_rd_en),
        .fifo_count(imu_count)
    );

    logic [511:0] lidar_interpolated;
    logic [3071:0] camera_interpolated;
    logic [127:0] radar_interpolated;
    logic [63:0] imu_interpolated;
    
    logic lidar_valid, camera_valid, radar_valid, imu_valid;
    logic lidar_interp_error, camera_interp_error, radar_interp_error, imu_interp_error;

    interpolation_calculator #(
        .DATA_WIDTH(512)
    ) lidar_interpolator (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .packet1(lidar_packet1),
        .packet2(lidar_packet2),
        .start(lidar_matcher_done && !lidar_matcher_error),
        .interpolated_data(lidar_interpolated),
        .valid(lidar_valid),
        .error(lidar_interp_error)
    );

    interpolation_calculator #(
        .DATA_WIDTH(3072)
    ) camera_interpolator (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .packet1(camera_packet1),
        .packet2(camera_packet2),
        .start(camera_matcher_done && !camera_matcher_error),
        .interpolated_data(camera_interpolated),
        .valid(camera_valid),
        .error(camera_interp_error)
    );

    interpolation_calculator #(
        .DATA_WIDTH(128)
    ) radar_interpolator (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .packet1(radar_packet1),
        .packet2(radar_packet2),
        .start(radar_matcher_done && !radar_matcher_error),
        .interpolated_data(radar_interpolated),
        .valid(radar_valid),
        .error(radar_interp_error)
    );

    interpolation_calculator #(
        .DATA_WIDTH(64)
    ) imu_interpolator (
        .clk(clk),
        .rst_n(rst_n),
        .t_common(t_common),
        .packet1(imu_packet1),
        .packet2(imu_packet2),
        .start(imu_matcher_done && !imu_matcher_error),
        .interpolated_data(imu_interpolated),
        .valid(imu_valid),
        .error(imu_interp_error)
    );

    data_assembler assembler (
        .lidar_data(lidar_interpolated),
        .lidar_valid(lidar_valid),
        .camera_data(camera_interpolated),
        .camera_valid(camera_valid),
        .radar_data(radar_interpolated),
        .radar_valid(radar_valid),
        .imu_data(imu_interpolated),
        .imu_valid(imu_valid),
        .fused_data(fused_data),
        .valid(valid)
    );

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            error <= 0;
        end else begin
            error <= lidar_matcher_error | camera_matcher_error | radar_matcher_error | imu_matcher_error |
                     lidar_interp_error | camera_interp_error | radar_interp_error | imu_interp_error;
        end
    end
endmodule





